//Udhav Varma (211120) and Shubham Anand (211020)
`timescale 1ns/1ps

module InstructMem (rst , clk , read_addr , write_addr , write_en , data_in , data_out);
input wire rst, clk, write_en;
input wire[31:0] read_addr, write_addr, data_in;
output wire[31:0] data_out;

reg[31:0] store [65535:0];

initial begin
store[0] = 32'b00000000100000001000000000100000;   
store[1] = 32'b00000000101000001000100000100000; 
store[2] = 32'b00100010001100101111111111111111;  
store[3] = 32'b01100010010000000000000000001101;  
store[4] = 32'b00000000000000001001100000100000; 
store[5] = 32'b01100010011100100000000000001001; 
store[6] = 32'b00000010000100110100000000100000; 
store[7] = 32'b10001101000101000000000000000000;  
store[8] = 32'b10001101000101010000000000000001;   
store[9] = 32'b01111010100101010000000000000011;   
store[10] = 32'b10101101000101000000000000000001;   
store[11] = 32'b10101101000101010000000000000000;   
store[12] = 32'b00100010011100110000000000000001;   
store[13] = 32'b00001000000000000000000000000101;   
store[14] = 32'b00100010010100101111111111111111;   
store[15] = 32'b00001000000000000000000000000011;   
store[16] = 32'b01100000000000000000000000000000; 
end

assign data_out = store[read_addr[15:0]];

always@(posedge clk) begin
if (write_en) begin
store[write_addr[15:0]] = data_in;
end
end
endmodule